//*********************************//
// 3p Vending Machine Testbench    //
// Jeph Mari M. Daligdig           //
//								           //
//**********************************/

`timescale 1ns/1ps
module vendo_3p_tb();

reg rst;
reg clk;
reg p1;
reg p5;

wire disp;
wire change;
wire [2:0] cstate;

initial
begin
	clk = 1'b0;
	rst = 1'b0;
	p5 =1'b0;
#20 rst = 1'b1;
#20 rst = 1'b0;
#20 p1 = 1'b0;
#20 p1 = 1'b1;
#40 p1 = 1'b0;
	 p5 = 1'b1;
#20 p5 = 1'b0;
#200 rst = 1'b1;
#20 rst = 1'b0;
#20 p1 = 1'b0;
#20 p1 = 1'b1;
#20 p1 = 1'b0;
	 p5 = 1'b1;
#20 p5 = 1'b0;
#200 rst = 1'b1;
#20 rst = 1'b0;
#20 p1 = 1'b1;
#60 p1 = 1'b0;
#100 rst = 1'b1;
#20 rst = 1'b0;
#30 p5 = 1'b1;
#20 p5 = 1'b0;
#100 rst = 1'b1;
#20 rst = 1'b0;
#20 $finish;
end

always #10 clk = ~clk;

//Main Code Instantiation
vendo_3p dut(.clk(clk),
			.rst(rst),
			.p1(p1),
			.p5(p5),
			.disp(disp),
			.change(change),
			.cstate(cstate));
endmodule

